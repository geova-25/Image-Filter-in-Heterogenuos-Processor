// interconexion.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module interconexion (
		input  wire        clk_clk,                          //                       clk.clk
		input  wire        hps_h2f_mpu_events_eventi,        //        hps_h2f_mpu_events.eventi
		output wire        hps_h2f_mpu_events_evento,        //                          .evento
		output wire [1:0]  hps_h2f_mpu_events_standbywfe,    //                          .standbywfe
		output wire [1:0]  hps_h2f_mpu_events_standbywfi,    //                          .standbywfi
		output wire [12:0] memory_mem_a,                     //                    memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //                          .mem_ba
		output wire        memory_mem_ck,                    //                          .mem_ck
		output wire        memory_mem_ck_n,                  //                          .mem_ck_n
		output wire        memory_mem_cke,                   //                          .mem_cke
		output wire        memory_mem_cs_n,                  //                          .mem_cs_n
		output wire        memory_mem_ras_n,                 //                          .mem_ras_n
		output wire        memory_mem_cas_n,                 //                          .mem_cas_n
		output wire        memory_mem_we_n,                  //                          .mem_we_n
		output wire        memory_mem_reset_n,               //                          .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                    //                          .mem_dq
		inout  wire        memory_mem_dqs,                   //                          .mem_dqs
		inout  wire        memory_mem_dqs_n,                 //                          .mem_dqs_n
		output wire        memory_mem_odt,                   //                          .mem_odt
		output wire        memory_mem_dm,                    //                          .mem_dm
		input  wire        memory_oct_rzqin,                 //                          .oct_rzqin
		output wire [7:0]  pio_0_external_connection_export, // pio_0_external_connection.export
		input  wire        reset_reset_n,                    //                     reset.reset_n
		output wire [11:0] sdram_wire_addr,                  //                sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                    //                          .ba
		output wire        sdram_wire_cas_n,                 //                          .cas_n
		output wire        sdram_wire_cke,                   //                          .cke
		output wire        sdram_wire_cs_n,                  //                          .cs_n
		inout  wire [31:0] sdram_wire_dq,                    //                          .dq
		output wire [3:0]  sdram_wire_dqm,                   //                          .dqm
		output wire        sdram_wire_ras_n,                 //                          .ras_n
		output wire        sdram_wire_we_n                   //                          .we_n
	);

	wire  [31:0] nios_data_master_readdata;                                   // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                                // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                                // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [24:0] nios_data_master_address;                                    // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                                 // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                       // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_write;                                      // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                                  // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                            // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                         // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [24:0] nios_instruction_master_address;                             // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                                // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire   [1:0] hps_h2f_axi_master_awburst;                                  // hps:h2f_AWBURST -> mm_interconnect_0:hps_h2f_axi_master_awburst
	wire   [3:0] hps_h2f_axi_master_arlen;                                    // hps:h2f_ARLEN -> mm_interconnect_0:hps_h2f_axi_master_arlen
	wire   [7:0] hps_h2f_axi_master_wstrb;                                    // hps:h2f_WSTRB -> mm_interconnect_0:hps_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_wready;                                   // mm_interconnect_0:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	wire  [11:0] hps_h2f_axi_master_rid;                                      // mm_interconnect_0:hps_h2f_axi_master_rid -> hps:h2f_RID
	wire         hps_h2f_axi_master_rready;                                   // hps:h2f_RREADY -> mm_interconnect_0:hps_h2f_axi_master_rready
	wire   [3:0] hps_h2f_axi_master_awlen;                                    // hps:h2f_AWLEN -> mm_interconnect_0:hps_h2f_axi_master_awlen
	wire  [11:0] hps_h2f_axi_master_wid;                                      // hps:h2f_WID -> mm_interconnect_0:hps_h2f_axi_master_wid
	wire   [3:0] hps_h2f_axi_master_arcache;                                  // hps:h2f_ARCACHE -> mm_interconnect_0:hps_h2f_axi_master_arcache
	wire         hps_h2f_axi_master_wvalid;                                   // hps:h2f_WVALID -> mm_interconnect_0:hps_h2f_axi_master_wvalid
	wire  [29:0] hps_h2f_axi_master_araddr;                                   // hps:h2f_ARADDR -> mm_interconnect_0:hps_h2f_axi_master_araddr
	wire   [2:0] hps_h2f_axi_master_arprot;                                   // hps:h2f_ARPROT -> mm_interconnect_0:hps_h2f_axi_master_arprot
	wire   [2:0] hps_h2f_axi_master_awprot;                                   // hps:h2f_AWPROT -> mm_interconnect_0:hps_h2f_axi_master_awprot
	wire  [63:0] hps_h2f_axi_master_wdata;                                    // hps:h2f_WDATA -> mm_interconnect_0:hps_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_arvalid;                                  // hps:h2f_ARVALID -> mm_interconnect_0:hps_h2f_axi_master_arvalid
	wire   [3:0] hps_h2f_axi_master_awcache;                                  // hps:h2f_AWCACHE -> mm_interconnect_0:hps_h2f_axi_master_awcache
	wire  [11:0] hps_h2f_axi_master_arid;                                     // hps:h2f_ARID -> mm_interconnect_0:hps_h2f_axi_master_arid
	wire   [1:0] hps_h2f_axi_master_arlock;                                   // hps:h2f_ARLOCK -> mm_interconnect_0:hps_h2f_axi_master_arlock
	wire   [1:0] hps_h2f_axi_master_awlock;                                   // hps:h2f_AWLOCK -> mm_interconnect_0:hps_h2f_axi_master_awlock
	wire  [29:0] hps_h2f_axi_master_awaddr;                                   // hps:h2f_AWADDR -> mm_interconnect_0:hps_h2f_axi_master_awaddr
	wire   [1:0] hps_h2f_axi_master_bresp;                                    // mm_interconnect_0:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	wire         hps_h2f_axi_master_arready;                                  // mm_interconnect_0:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	wire  [63:0] hps_h2f_axi_master_rdata;                                    // mm_interconnect_0:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	wire         hps_h2f_axi_master_awready;                                  // mm_interconnect_0:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	wire   [1:0] hps_h2f_axi_master_arburst;                                  // hps:h2f_ARBURST -> mm_interconnect_0:hps_h2f_axi_master_arburst
	wire   [2:0] hps_h2f_axi_master_arsize;                                   // hps:h2f_ARSIZE -> mm_interconnect_0:hps_h2f_axi_master_arsize
	wire         hps_h2f_axi_master_bready;                                   // hps:h2f_BREADY -> mm_interconnect_0:hps_h2f_axi_master_bready
	wire         hps_h2f_axi_master_rlast;                                    // mm_interconnect_0:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	wire         hps_h2f_axi_master_wlast;                                    // hps:h2f_WLAST -> mm_interconnect_0:hps_h2f_axi_master_wlast
	wire   [1:0] hps_h2f_axi_master_rresp;                                    // mm_interconnect_0:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	wire  [11:0] hps_h2f_axi_master_awid;                                     // hps:h2f_AWID -> mm_interconnect_0:hps_h2f_axi_master_awid
	wire  [11:0] hps_h2f_axi_master_bid;                                      // mm_interconnect_0:hps_h2f_axi_master_bid -> hps:h2f_BID
	wire         hps_h2f_axi_master_bvalid;                                   // mm_interconnect_0:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	wire   [2:0] hps_h2f_axi_master_awsize;                                   // hps:h2f_AWSIZE -> mm_interconnect_0:hps_h2f_axi_master_awsize
	wire         hps_h2f_axi_master_awvalid;                                  // hps:h2f_AWVALID -> mm_interconnect_0:hps_h2f_axi_master_awvalid
	wire         hps_h2f_axi_master_rvalid;                                   // mm_interconnect_0:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;             // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;          // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;          // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;              // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;                 // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;           // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;                // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;            // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_pio_0_s1_chipselect;                       // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                         // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                          // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                            // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                        // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_irq_irq;                                                // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, pio_0:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                              // nios:debug_reset_request -> rst_controller:reset_in1
	wire         hps_h2f_reset_reset;                                         // hps:h2f_rst_n -> [rst_controller:reset_in2, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> mm_interconnect_0:hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	interconexion_hps #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps (
		.h2f_mpu_eventi     (hps_h2f_mpu_events_eventi),     //   h2f_mpu_events.eventi
		.h2f_mpu_evento     (hps_h2f_mpu_events_evento),     //                 .evento
		.h2f_mpu_standbywfe (hps_h2f_mpu_events_standbywfe), //                 .standbywfe
		.h2f_mpu_standbywfi (hps_h2f_mpu_events_standbywfi), //                 .standbywfi
		.mem_a              (memory_mem_a),                  //           memory.mem_a
		.mem_ba             (memory_mem_ba),                 //                 .mem_ba
		.mem_ck             (memory_mem_ck),                 //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),               //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),               //                 .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),              //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),              //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),               //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),            //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),                 //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),              //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                //                 .mem_odt
		.mem_dm             (memory_mem_dm),                 //                 .mem_dm
		.oct_rzqin          (memory_oct_rzqin),              //                 .oct_rzqin
		.h2f_rst_n          (hps_h2f_reset_reset),           //        h2f_reset.reset_n
		.f2h_sdram0_clk     (clk_clk),                       // f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR  (),                              //  f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN   (),                              //                 .arlen
		.f2h_sdram0_ARID    (),                              //                 .arid
		.f2h_sdram0_ARSIZE  (),                              //                 .arsize
		.f2h_sdram0_ARBURST (),                              //                 .arburst
		.f2h_sdram0_ARLOCK  (),                              //                 .arlock
		.f2h_sdram0_ARPROT  (),                              //                 .arprot
		.f2h_sdram0_ARVALID (),                              //                 .arvalid
		.f2h_sdram0_ARCACHE (),                              //                 .arcache
		.f2h_sdram0_AWADDR  (),                              //                 .awaddr
		.f2h_sdram0_AWLEN   (),                              //                 .awlen
		.f2h_sdram0_AWID    (),                              //                 .awid
		.f2h_sdram0_AWSIZE  (),                              //                 .awsize
		.f2h_sdram0_AWBURST (),                              //                 .awburst
		.f2h_sdram0_AWLOCK  (),                              //                 .awlock
		.f2h_sdram0_AWPROT  (),                              //                 .awprot
		.f2h_sdram0_AWVALID (),                              //                 .awvalid
		.f2h_sdram0_AWCACHE (),                              //                 .awcache
		.f2h_sdram0_BRESP   (),                              //                 .bresp
		.f2h_sdram0_BID     (),                              //                 .bid
		.f2h_sdram0_BVALID  (),                              //                 .bvalid
		.f2h_sdram0_BREADY  (),                              //                 .bready
		.f2h_sdram0_ARREADY (),                              //                 .arready
		.f2h_sdram0_AWREADY (),                              //                 .awready
		.f2h_sdram0_RREADY  (),                              //                 .rready
		.f2h_sdram0_RDATA   (),                              //                 .rdata
		.f2h_sdram0_RRESP   (),                              //                 .rresp
		.f2h_sdram0_RLAST   (),                              //                 .rlast
		.f2h_sdram0_RID     (),                              //                 .rid
		.f2h_sdram0_RVALID  (),                              //                 .rvalid
		.f2h_sdram0_WLAST   (),                              //                 .wlast
		.f2h_sdram0_WVALID  (),                              //                 .wvalid
		.f2h_sdram0_WDATA   (),                              //                 .wdata
		.f2h_sdram0_WSTRB   (),                              //                 .wstrb
		.f2h_sdram0_WREADY  (),                              //                 .wready
		.f2h_sdram0_WID     (),                              //                 .wid
		.h2f_axi_clk        (clk_clk),                       //    h2f_axi_clock.clk
		.h2f_AWID           (hps_h2f_axi_master_awid),       //   h2f_axi_master.awid
		.h2f_AWADDR         (hps_h2f_axi_master_awaddr),     //                 .awaddr
		.h2f_AWLEN          (hps_h2f_axi_master_awlen),      //                 .awlen
		.h2f_AWSIZE         (hps_h2f_axi_master_awsize),     //                 .awsize
		.h2f_AWBURST        (hps_h2f_axi_master_awburst),    //                 .awburst
		.h2f_AWLOCK         (hps_h2f_axi_master_awlock),     //                 .awlock
		.h2f_AWCACHE        (hps_h2f_axi_master_awcache),    //                 .awcache
		.h2f_AWPROT         (hps_h2f_axi_master_awprot),     //                 .awprot
		.h2f_AWVALID        (hps_h2f_axi_master_awvalid),    //                 .awvalid
		.h2f_AWREADY        (hps_h2f_axi_master_awready),    //                 .awready
		.h2f_WID            (hps_h2f_axi_master_wid),        //                 .wid
		.h2f_WDATA          (hps_h2f_axi_master_wdata),      //                 .wdata
		.h2f_WSTRB          (hps_h2f_axi_master_wstrb),      //                 .wstrb
		.h2f_WLAST          (hps_h2f_axi_master_wlast),      //                 .wlast
		.h2f_WVALID         (hps_h2f_axi_master_wvalid),     //                 .wvalid
		.h2f_WREADY         (hps_h2f_axi_master_wready),     //                 .wready
		.h2f_BID            (hps_h2f_axi_master_bid),        //                 .bid
		.h2f_BRESP          (hps_h2f_axi_master_bresp),      //                 .bresp
		.h2f_BVALID         (hps_h2f_axi_master_bvalid),     //                 .bvalid
		.h2f_BREADY         (hps_h2f_axi_master_bready),     //                 .bready
		.h2f_ARID           (hps_h2f_axi_master_arid),       //                 .arid
		.h2f_ARADDR         (hps_h2f_axi_master_araddr),     //                 .araddr
		.h2f_ARLEN          (hps_h2f_axi_master_arlen),      //                 .arlen
		.h2f_ARSIZE         (hps_h2f_axi_master_arsize),     //                 .arsize
		.h2f_ARBURST        (hps_h2f_axi_master_arburst),    //                 .arburst
		.h2f_ARLOCK         (hps_h2f_axi_master_arlock),     //                 .arlock
		.h2f_ARCACHE        (hps_h2f_axi_master_arcache),    //                 .arcache
		.h2f_ARPROT         (hps_h2f_axi_master_arprot),     //                 .arprot
		.h2f_ARVALID        (hps_h2f_axi_master_arvalid),    //                 .arvalid
		.h2f_ARREADY        (hps_h2f_axi_master_arready),    //                 .arready
		.h2f_RID            (hps_h2f_axi_master_rid),        //                 .rid
		.h2f_RDATA          (hps_h2f_axi_master_rdata),      //                 .rdata
		.h2f_RRESP          (hps_h2f_axi_master_rresp),      //                 .rresp
		.h2f_RLAST          (hps_h2f_axi_master_rlast),      //                 .rlast
		.h2f_RVALID         (hps_h2f_axi_master_rvalid),     //                 .rvalid
		.h2f_RREADY         (hps_h2f_axi_master_rready)      //                 .rready
	);

	interconexion_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	interconexion_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	interconexion_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)       // external_connection.export
	);

	interconexion_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	interconexion_mm_interconnect_0 mm_interconnect_0 (
		.hps_h2f_axi_master_awid                                        (hps_h2f_axi_master_awid),                                     //                                       hps_h2f_axi_master.awid
		.hps_h2f_axi_master_awaddr                                      (hps_h2f_axi_master_awaddr),                                   //                                                         .awaddr
		.hps_h2f_axi_master_awlen                                       (hps_h2f_axi_master_awlen),                                    //                                                         .awlen
		.hps_h2f_axi_master_awsize                                      (hps_h2f_axi_master_awsize),                                   //                                                         .awsize
		.hps_h2f_axi_master_awburst                                     (hps_h2f_axi_master_awburst),                                  //                                                         .awburst
		.hps_h2f_axi_master_awlock                                      (hps_h2f_axi_master_awlock),                                   //                                                         .awlock
		.hps_h2f_axi_master_awcache                                     (hps_h2f_axi_master_awcache),                                  //                                                         .awcache
		.hps_h2f_axi_master_awprot                                      (hps_h2f_axi_master_awprot),                                   //                                                         .awprot
		.hps_h2f_axi_master_awvalid                                     (hps_h2f_axi_master_awvalid),                                  //                                                         .awvalid
		.hps_h2f_axi_master_awready                                     (hps_h2f_axi_master_awready),                                  //                                                         .awready
		.hps_h2f_axi_master_wid                                         (hps_h2f_axi_master_wid),                                      //                                                         .wid
		.hps_h2f_axi_master_wdata                                       (hps_h2f_axi_master_wdata),                                    //                                                         .wdata
		.hps_h2f_axi_master_wstrb                                       (hps_h2f_axi_master_wstrb),                                    //                                                         .wstrb
		.hps_h2f_axi_master_wlast                                       (hps_h2f_axi_master_wlast),                                    //                                                         .wlast
		.hps_h2f_axi_master_wvalid                                      (hps_h2f_axi_master_wvalid),                                   //                                                         .wvalid
		.hps_h2f_axi_master_wready                                      (hps_h2f_axi_master_wready),                                   //                                                         .wready
		.hps_h2f_axi_master_bid                                         (hps_h2f_axi_master_bid),                                      //                                                         .bid
		.hps_h2f_axi_master_bresp                                       (hps_h2f_axi_master_bresp),                                    //                                                         .bresp
		.hps_h2f_axi_master_bvalid                                      (hps_h2f_axi_master_bvalid),                                   //                                                         .bvalid
		.hps_h2f_axi_master_bready                                      (hps_h2f_axi_master_bready),                                   //                                                         .bready
		.hps_h2f_axi_master_arid                                        (hps_h2f_axi_master_arid),                                     //                                                         .arid
		.hps_h2f_axi_master_araddr                                      (hps_h2f_axi_master_araddr),                                   //                                                         .araddr
		.hps_h2f_axi_master_arlen                                       (hps_h2f_axi_master_arlen),                                    //                                                         .arlen
		.hps_h2f_axi_master_arsize                                      (hps_h2f_axi_master_arsize),                                   //                                                         .arsize
		.hps_h2f_axi_master_arburst                                     (hps_h2f_axi_master_arburst),                                  //                                                         .arburst
		.hps_h2f_axi_master_arlock                                      (hps_h2f_axi_master_arlock),                                   //                                                         .arlock
		.hps_h2f_axi_master_arcache                                     (hps_h2f_axi_master_arcache),                                  //                                                         .arcache
		.hps_h2f_axi_master_arprot                                      (hps_h2f_axi_master_arprot),                                   //                                                         .arprot
		.hps_h2f_axi_master_arvalid                                     (hps_h2f_axi_master_arvalid),                                  //                                                         .arvalid
		.hps_h2f_axi_master_arready                                     (hps_h2f_axi_master_arready),                                  //                                                         .arready
		.hps_h2f_axi_master_rid                                         (hps_h2f_axi_master_rid),                                      //                                                         .rid
		.hps_h2f_axi_master_rdata                                       (hps_h2f_axi_master_rdata),                                    //                                                         .rdata
		.hps_h2f_axi_master_rresp                                       (hps_h2f_axi_master_rresp),                                    //                                                         .rresp
		.hps_h2f_axi_master_rlast                                       (hps_h2f_axi_master_rlast),                                    //                                                         .rlast
		.hps_h2f_axi_master_rvalid                                      (hps_h2f_axi_master_rvalid),                                   //                                                         .rvalid
		.hps_h2f_axi_master_rready                                      (hps_h2f_axi_master_rready),                                   //                                                         .rready
		.clk_0_clk_clk                                                  (clk_clk),                                                     //                                                clk_0_clk.clk
		.hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.nios_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                              //                         nios_reset_reset_bridge_in_reset.reset
		.nios_data_master_address                                       (nios_data_master_address),                                    //                                         nios_data_master.address
		.nios_data_master_waitrequest                                   (nios_data_master_waitrequest),                                //                                                         .waitrequest
		.nios_data_master_byteenable                                    (nios_data_master_byteenable),                                 //                                                         .byteenable
		.nios_data_master_read                                          (nios_data_master_read),                                       //                                                         .read
		.nios_data_master_readdata                                      (nios_data_master_readdata),                                   //                                                         .readdata
		.nios_data_master_write                                         (nios_data_master_write),                                      //                                                         .write
		.nios_data_master_writedata                                     (nios_data_master_writedata),                                  //                                                         .writedata
		.nios_data_master_debugaccess                                   (nios_data_master_debugaccess),                                //                                                         .debugaccess
		.nios_instruction_master_address                                (nios_instruction_master_address),                             //                                  nios_instruction_master.address
		.nios_instruction_master_waitrequest                            (nios_instruction_master_waitrequest),                         //                                                         .waitrequest
		.nios_instruction_master_read                                   (nios_instruction_master_read),                                //                                                         .read
		.nios_instruction_master_readdata                               (nios_instruction_master_readdata),                            //                                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                         .write
		.jtag_uart_0_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                         .chipselect
		.nios_debug_mem_slave_address                                   (mm_interconnect_0_nios_debug_mem_slave_address),              //                                     nios_debug_mem_slave.address
		.nios_debug_mem_slave_write                                     (mm_interconnect_0_nios_debug_mem_slave_write),                //                                                         .write
		.nios_debug_mem_slave_read                                      (mm_interconnect_0_nios_debug_mem_slave_read),                 //                                                         .read
		.nios_debug_mem_slave_readdata                                  (mm_interconnect_0_nios_debug_mem_slave_readdata),             //                                                         .readdata
		.nios_debug_mem_slave_writedata                                 (mm_interconnect_0_nios_debug_mem_slave_writedata),            //                                                         .writedata
		.nios_debug_mem_slave_byteenable                                (mm_interconnect_0_nios_debug_mem_slave_byteenable),           //                                                         .byteenable
		.nios_debug_mem_slave_waitrequest                               (mm_interconnect_0_nios_debug_mem_slave_waitrequest),          //                                                         .waitrequest
		.nios_debug_mem_slave_debugaccess                               (mm_interconnect_0_nios_debug_mem_slave_debugaccess),          //                                                         .debugaccess
		.pio_0_s1_address                                               (mm_interconnect_0_pio_0_s1_address),                          //                                                 pio_0_s1.address
		.pio_0_s1_write                                                 (mm_interconnect_0_pio_0_s1_write),                            //                                                         .write
		.pio_0_s1_readdata                                              (mm_interconnect_0_pio_0_s1_readdata),                         //                                                         .readdata
		.pio_0_s1_writedata                                             (mm_interconnect_0_pio_0_s1_writedata),                        //                                                         .writedata
		.pio_0_s1_chipselect                                            (mm_interconnect_0_pio_0_s1_chipselect),                       //                                                         .chipselect
		.sdram_s1_address                                               (mm_interconnect_0_sdram_s1_address),                          //                                                 sdram_s1.address
		.sdram_s1_write                                                 (mm_interconnect_0_sdram_s1_write),                            //                                                         .write
		.sdram_s1_read                                                  (mm_interconnect_0_sdram_s1_read),                             //                                                         .read
		.sdram_s1_readdata                                              (mm_interconnect_0_sdram_s1_readdata),                         //                                                         .readdata
		.sdram_s1_writedata                                             (mm_interconnect_0_sdram_s1_writedata),                        //                                                         .writedata
		.sdram_s1_byteenable                                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                                         .byteenable
		.sdram_s1_readdatavalid                                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                                         .readdatavalid
		.sdram_s1_waitrequest                                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                                         .waitrequest
		.sdram_s1_chipselect                                            (mm_interconnect_0_sdram_s1_chipselect)                        //                                                         .chipselect
	);

	interconexion_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.reset_in2      (~hps_h2f_reset_reset),               // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
